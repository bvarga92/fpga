`timescale 1ns / 1ps
module log(input[6:0] n, output reg[6:0] nlog);

  always@(*)
    case(n)
      7'b0000000: nlog<=7'b0000000;
      7'b0000001: nlog<=7'b0000000;
      7'b0000010: nlog<=7'b0010010;
      7'b0000011: nlog<=7'b0011100;
      7'b0000100: nlog<=7'b0100100;
      7'b0000101: nlog<=7'b0101010;
      7'b0000110: nlog<=7'b0101110;
      7'b0000111: nlog<=7'b0110011;
      7'b0001000: nlog<=7'b0110110;
      7'b0001001: nlog<=7'b0111001;
      7'b0001010: nlog<=7'b0111100;
      7'b0001011: nlog<=7'b0111110;
      7'b0001100: nlog<=7'b1000001;
      7'b0001101: nlog<=7'b1000011;
      7'b0001110: nlog<=7'b1000101;
      7'b0001111: nlog<=7'b1000110;
      7'b0010000: nlog<=7'b1001000;
      7'b0010001: nlog<=7'b1001010;
      7'b0010010: nlog<=7'b1001011;
      7'b0010011: nlog<=7'b1001101;
      7'b0010100: nlog<=7'b1001110;
      7'b0010101: nlog<=7'b1001111;
      7'b0010110: nlog<=7'b1010001;
      7'b0010111: nlog<=7'b1010010;
      7'b0011000: nlog<=7'b1010011;
      7'b0011001: nlog<=7'b1010100;
      7'b0011010: nlog<=7'b1010101;
      7'b0011011: nlog<=7'b1010110;
      7'b0011100: nlog<=7'b1010111;
      7'b0011101: nlog<=7'b1011000;
      7'b0011110: nlog<=7'b1011001;
      7'b0011111: nlog<=7'b1011010;
      7'b0100000: nlog<=7'b1011010;
      7'b0100001: nlog<=7'b1011011;
      7'b0100010: nlog<=7'b1011100;
      7'b0100011: nlog<=7'b1011101;
      7'b0100100: nlog<=7'b1011101;
      7'b0100101: nlog<=7'b1011110;
      7'b0100110: nlog<=7'b1011111;
      7'b0100111: nlog<=7'b1100000;
      7'b0101000: nlog<=7'b1100000;
      7'b0101001: nlog<=7'b1100001;
      7'b0101010: nlog<=7'b1100001;
      7'b0101011: nlog<=7'b1100010;
      7'b0101100: nlog<=7'b1100011;
      7'b0101101: nlog<=7'b1100011;
      7'b0101110: nlog<=7'b1100100;
      7'b0101111: nlog<=7'b1100100;
      7'b0110000: nlog<=7'b1100101;
      7'b0110001: nlog<=7'b1100110;
      7'b0110010: nlog<=7'b1100110;
      7'b0110011: nlog<=7'b1100111;
      7'b0110100: nlog<=7'b1100111;
      7'b0110101: nlog<=7'b1101000;
      7'b0110110: nlog<=7'b1101000;
      7'b0110111: nlog<=7'b1101001;
      7'b0111000: nlog<=7'b1101001;
      7'b0111001: nlog<=7'b1101001;
      7'b0111010: nlog<=7'b1101010;
      7'b0111011: nlog<=7'b1101010;
      7'b0111100: nlog<=7'b1101011;
      7'b0111101: nlog<=7'b1101011;
      7'b0111110: nlog<=7'b1101100;
      7'b0111111: nlog<=7'b1101100;
      7'b1000000: nlog<=7'b1101101;
      7'b1000001: nlog<=7'b1101101;
      7'b1000010: nlog<=7'b1101101;
      7'b1000011: nlog<=7'b1101110;
      7'b1000100: nlog<=7'b1101110;
      7'b1000101: nlog<=7'b1101111;
      7'b1000110: nlog<=7'b1101111;
      7'b1000111: nlog<=7'b1101111;
      7'b1001000: nlog<=7'b1110000;
      7'b1001001: nlog<=7'b1110000;
      7'b1001010: nlog<=7'b1110000;
      7'b1001011: nlog<=7'b1110001;
      7'b1001100: nlog<=7'b1110001;
      7'b1001101: nlog<=7'b1110001;
      7'b1001110: nlog<=7'b1110010;
      7'b1001111: nlog<=7'b1110010;
      7'b1010000: nlog<=7'b1110010;
      7'b1010001: nlog<=7'b1110011;
      7'b1010010: nlog<=7'b1110011;
      7'b1010011: nlog<=7'b1110011;
      7'b1010100: nlog<=7'b1110100;
      7'b1010101: nlog<=7'b1110100;
      7'b1010110: nlog<=7'b1110100;
      7'b1010111: nlog<=7'b1110101;
      7'b1011000: nlog<=7'b1110101;
      7'b1011001: nlog<=7'b1110101;
      7'b1011010: nlog<=7'b1110101;
      7'b1011011: nlog<=7'b1110110;
      7'b1011100: nlog<=7'b1110110;
      7'b1011101: nlog<=7'b1110110;
      7'b1011110: nlog<=7'b1110111;
      7'b1011111: nlog<=7'b1110111;
      7'b1100000: nlog<=7'b1110111;
      7'b1100001: nlog<=7'b1110111;
      7'b1100010: nlog<=7'b1111000;
      7'b1100011: nlog<=7'b1111000;
      7'b1100100: nlog<=7'b1111000;
      7'b1100101: nlog<=7'b1111000;
      7'b1100110: nlog<=7'b1111001;
      7'b1100111: nlog<=7'b1111001;
      7'b1101000: nlog<=7'b1111001;
      7'b1101001: nlog<=7'b1111010;
      7'b1101010: nlog<=7'b1111010;
      7'b1101011: nlog<=7'b1111010;
      7'b1101100: nlog<=7'b1111010;
      7'b1101101: nlog<=7'b1111010;
      7'b1101110: nlog<=7'b1111011;
      7'b1101111: nlog<=7'b1111011;
      7'b1110000: nlog<=7'b1111011;
      7'b1110001: nlog<=7'b1111011;
      7'b1110010: nlog<=7'b1111100;
      7'b1110011: nlog<=7'b1111100;
      7'b1110100: nlog<=7'b1111100;
      7'b1110101: nlog<=7'b1111100;
      7'b1110110: nlog<=7'b1111101;
      7'b1110111: nlog<=7'b1111101;
      7'b1111000: nlog<=7'b1111101;
      7'b1111001: nlog<=7'b1111101;
      7'b1111010: nlog<=7'b1111101;
      7'b1111011: nlog<=7'b1111110;
      7'b1111100: nlog<=7'b1111110;
      7'b1111101: nlog<=7'b1111110;
      7'b1111110: nlog<=7'b1111110;
      7'b1111111: nlog<=7'b1111111;
    endcase

endmodule
