module add(
	input [3:0] in1,
	input [3:0] in2,
	output[4:0] out //out=in1+in2
);

	assign out=in1+in2;

endmodule
